`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VL5XljV1WG0oNRTZAe9MPv2ZybZ60ySrXyMSUIPAHCKNWHP6iO+/INtyBcE0RuzocdqTFG7sDgi0
VgofHyHOVQ==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
astDErvPrFoemv50z9CmdmoWPW5CNEC7bPLyuzZp6DXZsN98NXCm5toxXadFPVQpREiL5q7Zs7CR
BYsEz5B5MABJFUJCYxw8gisLp/RjHVqy4rUzLSSuxctPeeomal5hSlQh6POSXrzYFAo04FXxr0y1
/A3BDo7MBKj+MWXO2m4=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wY68/DQXKqyKNGg0Pj8ZlmPga7LglN+inyeDJzAsgOVCzxZtluWcygkpY6az0PRTvEifFvtJYY/o
BUzE2KGd6IIR6w1Bzrf49t/s5DSF1jALpSGCn0y0k2PLxcfsIYyEVlZLQAb5ycbEX3U/Ga6ikqBS
j63dRUfd9hCZVwn+ie1Ik/0o8bU4mIKdOeuwnEWzz53TJjjI16dPk1FYX5bOiRgHGWdq8VyInFkV
JyecGPLXVPlhlqJKjHKT4gcVZknBSunk91tx9RWaG6E+dMp4qZVuEQcVaB+yiDMZeaZkHDSsgjLS
c1EUeP2KE7Kim8RblcMAokD6HrfKuQHyMJIoxg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
i4ME/1/aXpUxAxwwPkLNu3Z9//ZhjvDRFPKctD3WJFh6t1WiSRmypW69atAGM6+7eldzTl/M8FgW
tx1kQwlIvRzWygW2r8hv9Pa/towQQ+QcvaY87c1eFr9NqzHQuizNT5hAM4toZO606BRXMasRn4x8
ZObqteLRCHL0H8XV/9KKfXxupyUqJyuYwfCAZoOxu0C5D806uA8vUjxQRzpAEBmR0zsO3RNOhznT
eVlA7cftNEE5fNgulENkRU2xmpKJt4kaxrVYiXKklzJ9y0x2jOxitzBwY/RHtQlysuVEGt769j+Y
iDR8PnPELFavy2DNa++LLNI7xlTtq8Gn0PHr7A==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jIySNDzqqNkGWmvkqbnuMKRVsQgwOzeVgAsWAHDPqDLFp2OHkwrgzsVw5x5sunJKSz2WffI9cZ1/
r1TtrI7HKxPplMfl15offG7GTfIazGLwHSEYg/X1pI+NwXdm1Y7V1JtZLtK7kaH3tngDy5+dTS7N
xA1wFc5mXgjeOO0kQa0PzDE8S6IPc6mXq58fJdm28SUP4dT8CD9+hw6+6N0EzOKBIkdBBYu8YERr
dYxUDCa9idwqRp2MlGcCkwLKJMW80G9NJukiVoO5jj2uglkLnaifTZfCvmAJMdmlQE3wiLnYjAH6
/5tLW3tK1djBZakJWAADYDvGN1Gfoq41DE9kaA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
htfz1DTXH+8I1PZWPRx59WNYv3sC0LKJ6q101DPCxtu3kx16B0n9I/iU/XlZfH8YtyYvYJA6YKgr
e+avYUZgNkE2POJTucOn/xXfMWqdUEWCaJw2neVEIESBJxwtc+ovBHgohwfLG04THjke/xYCDPnW
LIw4ZTipduowNh6rv08=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fX8qp7VCXYU+LxFYppmO9d8I712uGBvizO5m/RxD9yZRj9IyiyY8QH/iB3dZWraK0stmwE57MutP
umhrveyrzy00CNdWqmes2++k1BabPW+SNA9gWvvqJkKYHbM+aSRSVvnYEKF2+3i6m1i7Mocu/lW3
pm2nYwyt4Q6A7dzHWApGXcT466MQecgHt/gqmri+fbtDRMaxAUhaLMLOBxSS/Ix6WWU4hHVS6M9e
+kPiMt9xvMVg5Doi/B1U7gnW8hgLJJ6tDtC1tr3hwooqPAgXYLRDylhMVNChxxv1I/x/EEJfcjBT
r8BBAPLaxMJ16yjhu2A9LtJu0PAqGFIQf58nQQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10640)
`protect data_block
fS/hXSieRFR10bDf8kusVF1mmHhioS3sOT9/38r+TuNwXhBYcKbvvuKbnfR4DcTPJ8h36EjrGnBO
NgmQli1QnCi5bmQ7Pjft8AxGHfNr771+IMQMSs3gjpHD+sk8GYiHF3qipVCkqt8D6xkztV0jXxZN
nQbHP38L26DnA9ZSEoZ8e+aOH15fYuBiE5JfqnmA5aLgbAw0hnWMsd4RycddQNlufxZFgKuw/0dF
BvldI6fv3zLDCtgTRm7tJW4PDyZQgWP1AI6sbtVo0nrc5rPHuSFK9HRo3x1kSDpeKtRSybdzwHLY
M+35e6W0vgQxftCoxGn8WOt25Ogd8xqHU0NzbS/70FemAktVku8x+/e2RYtucqmKNHuJHM3l4sYo
vIRkFem215/kpmwVXWAOgBtkzKBKs6ZUuhYDqQTRyZt4K/nsRHlaGE4UJ+ONEpgfS6iSfZXrNg9G
+JlPIIFLl+/+DhKEUdKk8SwdjhjPo0o+rH2WDjfNxBL9aG1y4sGmYSs+Eps7Q/Qcb32eS5XMGx3z
0/6L43UskZ6LF+hQnd4Oz+iCJLIEX+HJxmVn060tGXVDACXcK54rDRjUFe/ckfgvUrW+61F9wl8A
PMzkAE9ZJmK8zlamyCOMCtxD4NH0xcfVv1+Td8ERirMh9ytH0brhrc3VpaFUQuFZ6GIj1F73VjGs
ZGIKKCSzhaHktG3seo2TU6Xa1SmvJ2AX0pHRpHMp/33mo+j0FP4XlvlaXA+siH9WJe2XeQDDOJnC
fgwLwTYPxzDdmh+9hyvSUM9UC5YO6mHK2nDFlTM6MDda62/6G6gNuhxkStsUJyUZHeA9wPdq82la
/xPd2VdfDef0pFDRVDnqRprkslNQvGmFhec2YDcasvCo2c7B6d0PLOmDptNZCkLyDdr4DxoP/9rI
YVHYsI8pKQjJKwE7Qbvh7qNbRmNLfUqZCFyGxabkh63P/8ziajgx3gejTRk1QMvTKZlai1P60g02
SPtHiGfycOTCU5YqJpM+EoIKl8Cg0MTqApCAFfBCpJy+IaS0k32VGr7nfCmox3l4sQyqIemApLSP
ldinqEVm+8D9Sh1syq/MBNBxZku/O/4kFfEkMWwdMbvtK8qa7vIW9NySFsLWuUsVkwqLsIj0Ozla
+F6w+Ux+uy4OjR9zz1nFZi2bMGf4gafS3YnEnfAPpm6M1nYjgDgUgIuqaIeA0Ot8fwZxuKkuEb3D
2tCpM6P70rwY7m18vd6iHtxzBKOJu5jm8IEthg52PPTyA2fYkhZt57I8JyI7B60636da8smhCSOw
TaBvqdhuu2rQN8bdXFf6Qts397ik9PFnz7bV8ITM45vMfD0FhTgQ9zZJ2QcNC3ibcwUR+oKRwW3l
V9WFVkP6lF/PFImCkd/NEBLpDcda7PkH26FqKqR0IZRjUBhFJ98Xoty9w4Tl6Db87/N9lLVSJ/dD
j4FQ3DGcxrhV0NOqO8os+hiqW2EVn3JSHidAPpXAxqgdbdIXOzcvcfSs19Uu1oHVT1+oOSC8uAUk
7xGJVD86rMGc436CiWy/LxKqv5XyCGrJNagIegKIlNSYliPeTOWXRMWAvhxxPJZ+q3NyC/eOQ7ek
Xy5s7nJDks9lS+CnSiQ+aUPtnYdX97VWZTUXdGDnHtSXANUshpcpz4NQSucvno1bJumOJjYoebQs
0m4UGirYOaHyu2cuk6HLNBecXztiYI6onvLI3GYEbpegBAkyw61IGBfIuru9fpBSe9zuKDfFkj56
zy2B4LqztS26JOCw3kis+rxqHtmh4hC842CjHeAbaw5I2u4DYZvcFayHtfIsf4dAxzdZHvy/RTZa
v23H6NEr++hailIKQRaltd5vZ+b9wJBQeP4bPwb5JB6hXj+nyROhvRhguZjHkbdH31c1mzzblwWG
Z3hr0lWp7tCao4d8MTWEa0Nzka01WJ1TcdIANWkhO5+Ht/sTAdJSjrJj4BHETm9O+tkQyfW0RXCH
Bsv4xKzmuK/UNgdwLtvknEPN5diYYT19hpaKXa31exwjk6/3EKjOrRYZTQNbd6e0bxP4rEYxSEN8
Y1ewekjopT72vZxW8tV+vokwXLcMSLENWP3EnCLJq0OGjjDA3aB8um0mtltEmxnBaQikIo95FMIA
yxThFBdGK19dsIBRqdTdU+iCkv1pcNI2/IeU8d9d8ySkIB+w1IIR1ZHWVnUlIgczVN5XMIF8Dp6e
T0sz8irF6NxwG5M1RNXTOgs72wdwg+VSY0oWsUd19TPaxu32EUl7nHMF7TMKZBq5njTaQPzwgQg2
O0iT0G4tdFMztfYIDem8s5fQ1ugRNAYLhq4NZxW7FVqnbU3dPT/LjCW2Ngw4Hue7PKRyE89rvX5J
H9/s5KnfYJokqfabNK4ELO61gySbSLLjAUT/eS/ZmZ8dBJf+fgC/Hlnkrg/AfRABg409kMtuWZ5l
KZe4ey8SxqaiBxOiyiXZGNgaUKu9yS1KkCmYl5aSMLcWvirV0XlKQdvfoT5PGwmcslto4NmVP79s
J89l2hKk9G/ydW0AHotRztfv69PpSSOzoL7BMSGGhpeYElGq6KXTOPTTenvFpALdMO0mOcTraNFB
hs8VWiIdS/Jf6gXbZEx+7oYF67NTLWxePAmDN8fIuYwYZAqoeclAF+S3Iaf0pSiYspkIxXApBr+i
ZB9IXgUMBLBvTFKVXv6vcrGyKw0bhReMsOFk/ca0LDSyCjcpHQjdiwELUdrMTje9+7p3ziSFaS/+
SkFzbwsl3g6h+z9ORwXJSdc2rFrg4pAN8lNen4DcnJq5dnvo3ImPW0GeXSFF7ObkgMg791uRGocK
rd0+7r+UVVsU2GVko3Naq8Bc8BYZFcLgG4U+az59fAnusqNCl1WtbIDzgNvmRR4lcHnACLeh0yv5
WvSzm7LVuxRh89QGPiTBB7BHCIQlP24RjuOoeY+gCJQcLALvdecKQXRMnbnPF5TDPl413vUHCobM
CjIsOZzkvGaXpfIGDIu6TXdik+Rj56EvvWIew3ytRnLeq0DTEeYagGH+9fxBn41e+Fo2YMBJYJJI
cbmwA6pHoU7rx32h03gaFcmaRjF1wFRPtqsHyXZAFtsJcP3JN9Yl+bM8RVjvKlmTy09/1HOpOQZF
fNetW2StdbumRdGnTvJKGDrI3Fs6Iqz0mh84zCmeamNFZHOVbOhUIm6OTKsCZHmYvRZnzkepVmus
1nQq4vOe4iI9YypnIyHfN9AEBN6iMuarUgIoBmm5yxTZ59hrXG4gwggGXH0S8QdhKxoA+w5fUL4/
E1o3155tqyFjCMOUgfszn82Ck+jV7L5ZjQqiqXaMe9IiDiv1+dwcmE9FuP2UJfVEGZXKQTi2qIwd
/AkN41AXIW+3ahT2TE6W49DAjy/V/Vutcc/CuAlHSBdvGLiBT4NhK4UnebKWtkHRndvoOKN494du
FacdlbfeTqLFEfZJJ+ZFHxHYIrAR5KQ5tggz+8PxqW9PSTVM50kR02uDSvMA+/ZuGaffuBu/Rex8
XRBSIMqFPvBc9rArl7ydlXnQY9szeiKf5L9uSq4J1xNymbS9wpr3ucJXGJXMHlNrD1CE0P2K5qbg
h1hb/E5Esh0+ucr+eAKmyO1Uleyry8B25mmC8dhW2OgKglk1/2VrBuXyUdH0O4ArN9/LGmqtvvW0
NaDmwfIspivpl/PvzYQq3jaLfJ/nR7oBvInAJFrGQ9Sqml6X4nkYmXHJp32LzeGPJHRoimTgDb31
E2GJ5QDIrsJapN6FwvvQunGhLXh/fqtS8CBUjiTP8nh3UtmOPSkcBwGHU1kWHZOZ7JlHpD4dJKpQ
olbHhd/nTWEGwS4anGAdfaNSM7ae9WmuNCugMinNYN9buaAbNNG4S0xe0cjyN2/Qda2YVSnUS5Vo
ewmIpw2rseRjmDSu1IUWBACNWniOJGl9O0Q03vyZVMqpfyuZBnF8THGtMem+Gr0/CuDJyUeWKx2h
db53SgF19fkxo0FnfztNog9fU36tjXAQJ+ntGT29zkMnALq2H4YKd9pldRmEy31eTDr81NiIXzLr
uNzlnFdQnkjdXBdBftvLa0VM0cabD/hND8Raj6fSM64PAxV4sAeIuUKef6EMV78WMV8sc8OaVrTm
9kyW6+m734MMLa1RCvf3FnPh5J706WBL76fyxjmL1OlcDsky9CADn2TQb4T73w4tQ6+36eYldO01
j4VY7BLpYHoLp4yJgv3EZywxFU/aN6eU3e/O6fB12eeXXy5pcUgdMu0DLYaOadVudDRA0h4ktgMQ
Ngee5oqpMKvd8RKvWk+SfUgphbM3izEv2PrTVnN6Mioov0ARzBmZ0Z2VJYv7mY1xuQqj1Aog71Z7
wJegQdyIXa7nVJ1cH5aOTGDqt2pzVIxCm60h3tIB7obBhJRxXSc0cT0V/GodyHvaN0g97DZKZtaV
g7doEju6ZTR+Lq//0y/tedPdwjQAtzUGAHJs/0KHoCQBJ6RqNQLn7mJfpyU9liillp7w+SfhbnAl
T9mNQaCV9GlW1UW58C+hUSVXMd7FP/Z6dehlIwbJ3EyjPv1FXfl91ObJ8k+PrJBfa2V1FdGNV+Vp
e42t6i0dVEvPoeJ5q9ohIYC/iaI4c9HIifDFme+mq7LqOL69j1drlKRYni+nGYmAifJkpcUogk66
/mNuSYz8xTUSyZmTNOKB+Jggan+QNCaW21QUMhCazS4tjdvw9896WLV35u4iEZZ4fhVTHSyt8Cu8
6JhiCTLKWgmkB7IyjutOc4GuFLNV47E4dDneoBdGQ5IPyyalgIEKHliS9EbGsipekOuoxVaJJoQJ
KE7Dktgpf3YeK7XKt5kBox1pBL1TBXpOQZzKWEBHfbeCDblvIdb8Evf0Py+TiwMyimVRqrgE3B9d
ObNS14CQI5vxFQXGOHTQhNoh24FcHKACg/FykX35BfQ8dkq5Is+xOjTGYc4It/gVhPJVk02mGej1
Fs0w0XMcbWLXz2tGl+mCbPOUDEhd40IXNDd9rGq5TcpDwgwM1o3u45H+s0/9WYGUlDOGKrPoacnT
LVuRd8vNmPSYrCXcrFLdYveOdO+a0+uSyT+Cb7MzALeJSnkik5G2hTNS+DePeiRRrDvedtCY6nqg
1ns87OImWIFijGQb7sJswkzgH7U/y0ypH73YutZ8cOlZ18va8Vg4vZIqsSg1XdxoAB3mSkBAdYsF
i3w2+9C6nzp7ZU/E+PDMhUagPsfy/R4CH58KxgkcTPVjq+Un4fhX43nkfqQMNMrVFlq90Kmb1aWW
l1R5c7WS9tpi9EKuete7A5yjJJ4Sq1SFH1njvsgI/kGtgmQUG+5wxCuxI1Nc3KB7C6enlQBsmqKL
luHXyF65LAJSd+/0bi1A6OVNpKItcZnXRSzfTReZxskA9kkz+5EFMOtXQEr/zA1XXNzM+xBHktoc
mwKETXUbTfdzpzcnMFstQ3SzzfMvcJQ0UHTLPvnd8vSmMYC5yG2kEF/pmevjs1+p1mLX6L9EYW0Q
oArSw5sA6EynujdPf1NbmBS5fSXXYT3rFKCVsL15Qv25qmoEj+3pgpyzaYhDDBgc1qEJsznTkWCK
zptPY9cDX1KFb3V3ieycUJ8kOnQSK/z51d7AUKaBNntuq/dbPALipVO0i0IKnfP2ef6bNqOjx5mg
NAAH9jD9GQk8HAZ5C139mVVylxohXCYaHR0Sl3Axn07ED/1ChLOOQb0Y+Izbow3g0b8J8DNgarnK
qldgCGUqCWsx3Af6j6xsxUsqfMGsFhOa05O9EHvlLZpkYqpMvi0CyzPdDxM0TNQFHeocx4KfhqeZ
Gmcsf/hCK2kS66awKpoIZxxhVFo3LEB47JOh1M3cWIKX+0fSFMEZPKFjFK6Q6oJr+KnmRcMJE7lx
Q6zNDRdyVssOpb+RmAJNnbJzaxQ7LqHYPzhKm/mkFq314TPVAbWxmpGt4bh6+1E3NlO6ZW8+fdY8
B19nByzA1iJsYnAoNainDlzU819o043Xz10XIqvz0GBwqxJTxYMOtNc1v4i9+HiWN/uAjS8kS2mH
EDFWpkgKTSHnswbdI4KkHOQHzH+QhVMy1GOYABv5QinKsxFXybugXDklXrHqDZUP/Io7N3J0sud4
G2SRdwfNMwP4xxbGzSlhAGt2rnKEzY8I9DPhGp8ka1x7WcTxjdeXA7CPVWTMSjlPFHrgW7+JXNkn
+AHZfIbVI/uNyDKm0QgWaJPWKzxiIo/mDn0Vt46hX2UmDHkGKFpiRlK30XxFTRs5owTQeQ4RpKbB
k+FS/fl3GVsuu0PMDSPvTb6IbndR+RqfkVBp8zz9v4Bfc8A+tcPsKTOwZUZ/JIEeTC8PVRTu2fXs
+gD765cQkaB6Lj/YiwRsVyaUFu7DCwqH6lzX448Yk6zJ/PNr3iWdmxWzmArlV5n6lQVc0JLZlx6Y
ZaNMjzAK0gd2LbIVKrrI98JCxDu3/9iy1LQXhWSrREF2Db97apJjCRmbEx/8zNgKdycrM5eTjWln
MSrgtzg1xCp4XYxyrQE+PNrcqE0KXxhvW8z1qvSaiPU5tj313M89wCV4gz57elkf6WoATxtLOIzz
+bLHI9mIS0u4LOx+xpC2ENpZTR7hZ/UYdjCDE9o2v+4wVEwYK8WXzyPZVdrzF5ZV2fgt59w3W6F8
GZO+X8Ii7eAuYAkMF7psDSINDHi9uy1W8LnDC0EEfbv4BYLmPYvnWc6q8UKkWR/rWadTmaMaWdf7
tRX5MfFrJpplyFdHVS0EojkUVFIxm5OkvSmPwSXNxlQq8p32EaIXlGguftGo5A0dAa6gwjt9LdNb
EUYFto6RARrTpm1KGWP9MghBNYk09v6wfOmVTciH7mSC8oZGIr+nayBbCTdgrAnYwhT4WAzghNaV
NsLdctpuxodFohHcZsNHZpLfE4+rpdBDJi7IpUz//W50E9Gy8/wWl7tyv+C9M2kxKvtL+hq/1uNd
f5cJsygcjukmLMyF6qvI2dwtzFU+522qzxzZyJZh8PolafvUr3BjhoJYL7OXZz40VhtMWWIXl2JA
bVpM6fdJa7Pmj/57/aQeRPPLPKACUQLCDWZxdGbmC9mAP8ZUzMmJADj55D5fTMdj3syfxVyJyn8k
n+uGOoOs48dAd0lVYaS/A603DWVjMKsjCA9tZFd1u06eZ0Hb0bSPLvOZg/JnkI6hkthiP19PFzS7
ZMk8q7i6tvcdfxF++4hBUWJKzPnU6/F5+HbgjsRcJt59JUR/yqBzJ6N8guJyWdykyew+dZEBE0Cj
BEMPg/v5GDoawS9tUJUuBEWR/DA7rtlFeuVEyL7yo70afQhEtmzPFBboqD2neNSdTmkWVq/1MHqq
tCK2IUpPI96PBbWDDmvvHCDbF0gZGOZ0HeZHTnBfcVtZ8xF+MZTQbsm7MLu24k4ZzwBnOC3xzR2W
bQeybshMeD+XCi5O63JVZax6gpnH8mGw4VI2gNQfWsWJvajthbTbgl7EcNxUKWU6JKgSUb5ktKJB
iArCg54D802oY9ObVXGpPYa7tThHM7EbS0WZhnkuInFQakQ+m07bNKAwLkEr6iJXN9hIBIbz7pCW
9phTDdEZHsWJIVfMAR4XhobDyRe4T0EikRrpegC22ML4A9j7bxWm7mi0dePPCCKtq76uHn4gZm3I
BDtXo9M1WuzOFgGdJuMtv7evmG44e2uxS+AQ7U+uhRvma+3KU/B5NeknmS/0WhxPBkPiMxb5aP8Z
4gdggio8g9LUfng90CIpY36KeoKQeNb8mzlpgmPdsvBBDUgM364LWiuBLtHsk+s78lj0zrE/vxjh
MFu409BCPM6Yyt4M2UKR3olmLH/yz6Q3HKNrAp7sYFsxgu0s5Dy2YCc8tpiOiaJkFz3AVST1JqZz
/622Ms2qn2YgvF+1Zw/yILLXeBWyAIomoYzJ0I34RBTSjHyw3iMM9D9GL44MVv6MjrpDvxx7c3ci
xyylqE4x+7gpkQalyBAzogXYLTrV87+FdES2Dh3QydQf0sQW9ZwkqB0Ba9VD7bnR34ztyTiAdYIs
Ft9Jwpvj45EJRUHAqMNL3fnis1ElsNy+UFfqXBVXKuIeYm4UwaLawKfep7wfN8CJ0ScH4O2u1Eyp
zjlVVPvA7r+auzXudiwz9pNN96PLAX0ofn5DHM5MgF08az+nxdIGX+aaRNkHHFjr18RgltTNLuw6
uiKpK6AjY9RcvffR06fhQrlDEQesxpRBjtP2pMMUBaiD5kv7DtNhwBvofltU6a0D5PRonhIz7Oj0
rR1GJw7kT9xn3aAjgcRw78osVeyJ381COioJhvf94OIFl6i51M+VkaVum5maChrnfozFjGMBzfjZ
cS/6UlqPTcegWkr0gk5izpy0LPDuYb0V0LYsdvUKCEEFnDQENs0T+qLyjXn0i4otjXegl9QdIWSv
lYSN34Pjh8rU94rRe3G/A+O7RKJapYyAYRvVjDRrq2nPjKTr7Wtjd5fWT195z167VGLnMrmqgp7y
8+rRE1rXjdHIRGg/hDg5HxveMj99uCU4bEjbCuH/UmWR9aNu7XIyUqI2z9foYAJn3L5vRt7kuumP
7ddkOTxaYRk+nt0SN+/bD2PEClpTY2/ZNNjHGj3rv5XQsxey+q3NwKPo6pLUHzD4LcUn/5p5VI9D
cGze/XM7bjeiWI9hcSDmVg1oIaJa9V/8iXIb/JBa8GDxETDHdcSb6K9CAnhnIupn8kw9PHu2fTJy
oMedBwBm814ngAkORxc0fI/6hgBdBYo+BjY0L8gbQjswPs29nCH042Jvhv3G0875k6nvtqBOUZNo
OzJph1Rdm6h098nzA1+bqCR+puJF3Nqd6+YUsZs0j2VTQ0MHtMvH9ZQAJSJcRcH/a059tFSDDzSC
knxVsQygIrldg3eiLZZpVxOHBNzd5NGyDgQlBZbziC7czNn/s9Vp/hRUOovnvDI2DYLqhXKLxoWm
uNd+Boq9+6HWxSKMBQBVBMSxBApqcQDUC+UU7Ku9bBG5F/kMVokOch33A1DKTC+/X4hswA171IQ8
TH12X9M52E/w2kT8IK+gmb+1s7IOehre0Eva+JJewYx5ueMeSkLrWCibZvUWkmcwFwtV+8Di3j2b
wxtHkEBdRQ9Y3Fgi3ksP39lA0CQObYULCXhikUwdkTpgYDquIWeF2YiMb2nwdAa1TzjpawpijpCL
gaUSOxX+TFcA1IjaQUUR/kAaPw44qzrj/WNCiC61yzqUPr8iChv7Iqx/1/F1p73NJKulWvvafrG6
lyYb3aXhmLqQ6a4QheOlGBSHU9CdsAcG7qc5qIFK4jkmB2wg9Lz/MrLOg7nNA3MKr59Uz+qx9Bc9
uJVj6WEsPan1gvLTIiQMvaRNV6kH17aCON0K1A6ZZAkThDqWZCxfveURSXg2n+kcPHWlRVInz8IU
ANtNZDGmNQvH1YRLd4PuNw/MAY75OHNlWG4oAl83HO5Olo20O+UCLeDjs2zYgDBCEnYlrCzcNDvg
hTaSf5dECsVz1X6nHiRMMVFLNupRyDwAmrwH68/uVWGD13cmpB8I3PQYa35mzpgdFLbV3YcEauuF
Pgcx/4/IVkvXxeWoaj55PD/3HEFSriA4p4sdSdUn/y+FX0QZsCVn8wreXnXYGdGw7GzRT577ZJgu
xWzecxjwF2tpHwn5wwzBdQmcdDyBGioeInz3IC2EkCYg9yToHeLO4XSz6GNeRdrbTTrsXRCDd1g6
ahdAEWGF1gYdl+1jR74xkKgerRyWqD1XwIwmnsV5u9N6//js+7jZ5qF/ku/LJ4RWk7S1/tcJq0FO
lJBm5BtRJ/NlexBW3EBwCYSB7gYVfxlTfCPG/RIbUsncDm5NqSiY9FErJdFQ1qwzufijjpXZjEKA
BakcTwKC5VpX18FhwQNl902lFG+37DJCXkWue7QCODbcSelgavXqlDRzZSYRQf/FjFD6xq7xIwD6
67yI5uFwhJiOX7V2V3L6kNm8EC+A1X/BsdSe8Eo+MTYrFnuNdcgdwX/ucWnok4Ubm5dRfwJdz+19
XgoTRW0CyGP6BVQF2MUz2CU2MTeda8YNAEQ8/ubVA57l7118oVNdfY/MhlLRIO8Sp+O3cvV+jBDb
kee0vgkhw7VNwi9Huo7IdpnmhAoAGcKplG3W2gCdp804pf6BjQbdFPwO1SnkhXz9lU8Ue42P0/bN
jjJyGWaQPJYqEyWUfCD4U0f2ukc7c9yjRz9lFEHFrIBCbRnn1DxHTWc/+3w3brHRPnQ9zEcS0QCq
39gaLPrAc/FDhAhYLODLR5fE0CP+JcPkDWJsdOMWCwrapSKj9FOQ0MkpS4kPnnBh7jq/X7fiJcG0
mkKUv/IjwMzntmxSzvoQcrPPsK3eKDOeCtY6UnAF3GsGX9A8rCQ+YCkK9c6NySM6fmoDuw1Q4z2W
3KoJodNlVJAoQ0+07Q9Qlbwh5OUrN+9wi+WNiwHERAWZtLm2H729yYv34Rh5TyUqnA7vSuJuJEAo
mTTHIBto7W93/0Vt42sx0vp5LONxJc4V80Y+TLRv6PkVboYLRlLpv4abXBhUZ12nzMuqf18IK7sZ
VOZLunjNW+X1byzOQFAbkB7QQ1Decc2F8mOiXv9zJex/yhJXx+OimxM8qkOnpqDIpitnNKw8SQV7
jLk8pm13ZH6bOdyIhUAEq6dPHKm1rRqUbWdEB/we1jdXdhtoYWXDAxuALrAV/1AwGzoIZMiR+BDm
VSeERTEDsyNh+uWQ0R8xgRtc13oChGILpviPWvzG9sx0BqdAmdwpdRSsqqHWF+MNBBPpWYcRY75V
dE9YxO+ipY6cB4aiuAvPbfRg7p04xdngaI0bk7LnJ7A5coqGp/9dat79y1bzv+ZaIDexS3+uz8Z3
R6Kc6JCud+mCOLJnTewsbXoCDgrVMs1i1gNOrgyJTdIMhaCibzckqvDz6kjFTUTLBFTzJTKkPQZa
kULyrYwOmZhKyQbOxh7c/l7bvvurOLBaZ0xG4gQUpKU7SCH2IDP7f+T03+IuIobsduIZQRP5os0V
JQjEIrdZO3syhOYYYrTuWTCUFTiGxU6lJ5dhsZUDUPjoBh/clkWc+B8kOKzOGSW+6f1YA7tx71xR
CJ7qZVV0Heat7qUOxcu6IbV/OlX3injKJbLBGD0Wo3o2V+yCzDYC1zLtSHtXMXcMSqSZG10w/Sid
lHsUEl1x7qLdEHyWWIvqZZf/jfz9Lfy4nrldt6Cp7J+dVfIWObrFfBkIh/y6WJZdy+fO6lOTzSah
yHpvl9pYJzjXPu5JzV7gutQXbWp0ugWvOiGtCPrSn+kkrI5N09v4u99oWKTX3QgV4IYAqEmXo6Ie
qOh3yp0LngacEQV3/k1Gwgv8Np/+hI9e1NXILIDySE8dMDlIdY1yTTc8dGR9hKkVI4xyUTd9aoBO
yBTVsRwMAsBghi54alitUMmIalOKcj6t1USug2OgSuW7YNG17ISeo0DS3/LAy/kJunEME/LSRBkD
qelWSHTHEyvrYGh5xub02d30xynUzvVbEdOM68bD99E6rz/OTxJStCq06rPTxwtro2ek4menkg8o
i6/cHoRRRXoE2tWmpwNUzyTDRHEHmHZgC8xoMPVz8YUAjDnKDxHVnL28+2JHyzwNX2uC84kTZ7Aw
YHFkezbLi0LFSc0E5aR6+TY9rEuC9exXAHfLaiKtSti1e4DtCGfTXt1RjVu8WBj3svwhvBc2KVoE
yjHBe18VAFEqWGE8Wmc3giLNq9hHGPrttUPfeSePorCtXwHXXFM8YNwMcsIXPTzGgYRm014MKaUL
lCb0QFMSEf1WGNYz326m54KFus/kB96WeO1y9j/zjfDEUO2T5iI+ABycVbGGORqf1czUtCtyPHKR
8mxQy2KcC19dI9I/b7lQLQuCxyN9pphSz9oEw6/3+5G7xJErksRBBcNfBlIPN/R3rNw5NHQcvOl6
OKLbqovIDs5LpCLf5VWTTn/f8pPRmIGHTwD2h9fy1J4JKKU4ETfyKzTB/tsOHBXrqpb3B9i3lVjv
44gan/dTJ6VlCLzHBUnbCvNKlggLjHPKDBil3ul+hM8hAFJNDTaPqLBpJs22ZiPjKq332TMRdyPB
rheF+3MuZu049sbnjM6OKJZNL3n9Zth7YWFT2hw0NqL5e+4noz3vWBnct2vQCO3Lum6nGLQgH85X
9SyrAlhkp0etkvoB1bVW7+0il2m9h2ll5+xFUoS9UPXhzUba0Gtl27S4Tq6DBKzXZOeo3+vk6+jv
/X1i6vv9uiXJ785V0Ic+bjh27uTH8r+Y/rW8W2mktc51fL4CxJ/pXvKFJvCWjlvE/yn6yzgGapkl
Mh4RnoDJbEzyTc9X9Famh7lP3hQEOrp+zYSn3X19sdSh05CG/Ot8nRM7pK+qmjtSPLLXqKIy4PRz
NeF55MaguLBKE9I16OW1S83XsgBdzbAYuFLpFuxRAAN//HK7wd6xGH3f8Zo2SmMxsmGQ3gJ6mt02
s7jhIG8Nv9DCaHuyjvIrpm/dyD3HggzMByTJeC4mBLGE8KTKwar75VfskbMNwo2jgP/EV6iR2FkK
NwJUSMTbOAIK/+hLyyBXsKOZDmp5G+fGUiQGX+Lp6sNvOSbL8wjiTk20kSouiv1Zc8Of8jlHan/q
k7DNaIrcf/NrO5Z7Q9DRZgJ2TAa737B0f9B5t/Xy2JHZrIZEWBHpnQnoVVGlmF4P5NZ3CN4zx9LT
zzPeF+M/5927g91cVWzbMu4b/BHs0kKtzcdDfTPzkMB7/VYh0QERsCZT1hJ7DBraAqOIX37kjSw9
eruD/1WEx5Zn7Zg7AFiad6qcDI8V36BePSOUSicuxWQZDcfRkZfAARc5YWzBdGfETLo+CARi4VFx
xHyMh4Hy8xEI/nclSWw7m0XcWwK4zM0sGLJFR4G9ZyHyCGz+E0RS6BEM9IhvfDcRZlbEkvmmdLsi
fMB5ImYza9jtzjOhuzREn671GWEGNp6TN4aLrW23oVTxX1uD1zZzDjclZscAUfFm41ZeFRKtHD8n
34u1hvWBAzhX9g4RzRayNFosCujRHy5M7ppnXerKZB6UrnVI4feKPVJ1yryb/ZwG1q456o/gjqHZ
AFwU0eE0rq6GLS1gNxiy7enJI4yqaMDiwkfIDRh38p5Lhmcdrx3M2Ldfp0hxcURX8z96/U/myV29
NKxdVUno7udYJxr79vVuDHEn43XdO6Xkwhy5HMqwA9fPp7Yv35GrIO0hRbjD6WEYIwK8N3bpMr4Z
ss5tqe53z3cz8hz/SY2irf4p0d3tEYXJFh4W5H6qenja8daGjcRNNZuQ79sUm8pajYy6gGDduoW7
pIgEmo2d7Pe6sHodwOEKYpBmTKBcjnDiYzjitKCIC0YDLYAXtOPqDGHQVZdIpehdyXKNEH2RtcnD
fJ6Xzapq7PjBHnSmXKrzFlkFEjYl350/UcK5O15xpnVS8l8uMAU+V8yc47Jvb8xwy3UHuyRyfHzI
JdpajVikvIzJyfTvajG4sjV0A4OtQgnXBJdaLvKhx9S9m46+aqxhecvCU1wrUGWk9y1F3AE4bLIs
n15bZqoQ+8GxpR9i+0zMicpPsjJ+zxJ4+S91NbFof2Ke/c2BV3AqhzK2OHs+glbgZrSlWiNuRL5w
uBKxDDRTOgOObTe+oVh5lSAXvDqY2JQ5f4gHJjDFyjOeqVsF9nhsFqP4mbzCvX1RrqlXvBwY0jRo
sr0hP7s2XdxUNFDqm/86t62EfSLpvY/1ZDu82gjE6m64eUGsnxJnbYFp3scAOj8PiCnln6RJIgb4
N7E+MI5M1xLdwr1s5Byb0x2lUNUm+dvJo7Jo0KN4HBB7nTEkslJj+BP9AchXVmZjymWv+5bCRACh
v65BX6yotuYu5+il5I13p+Jke+gaM2daywfn2NmbfIeIzyq23qGlZFoPN2HdFdPz4inhbeUO+aUP
LAeSQYxwtAcMSiNrOydVxnO62jz+8E5bXTeFNdXJC/rIaXtQRbzBZw/ltdCN1arnLB3UTgSjANPQ
T9RaO6ClJ27MXxSizlSq3LVnfEQyCtg2A1DO/HFXHPLdejUmwk6tXQgt1dJKYUn6T6P0OTaTSsde
PCoc0IKVpH3cy6yrsdEemC5x+VMdievki/8lP6mTXGFXQTa81Pc0AR7+XLiTKo3BUDJyQfS+5tGq
jPSu3J/dIa1764CNHDzDW2ZL/M8ohPZSL1RRLVv07QfH7eXnDNt/qAZYQe80LEZWGqfl5JIAIKsd
DG1E8pdqLGNcKOavO/PJHCh2PIkjIk08Hd8CrbHBPJN0BF5BcgY=
`protect end_protected
